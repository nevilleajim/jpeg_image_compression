----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12/14/2025 02:18:41 PM
-- Design Name: 
-- Module Name: jpeg_type_pkg - rtl
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

package jpeg_type_pkg is
    subtype coeff_t is signed(15 downto 0);
    type block8x8 is array (0 to 7, 0 to 7) of coeff_t;
    type block64 is array (0 to 63) of coeff_t;
    
    type dc_code_type is record 
        code   : std_logic_vector(8 downto 0);
        length : integer range 0 to 9;
    end record;
    
    type dc_luma_array is array(0 to 11) of dc_code_type;
    constant DC_LUMA_HUFF  : dc_luma_array := (
        (code => "00",          length => 2),
        (code => "010",         length => 3),
        (code => "011",         length => 3),
        (code => "100",         length => 3),
        (code => "101",         length => 3),
        (code => "110",         length => 3),
        (code => "1110",        length => 4),
        (code => "11110",       length => 5),
        (code => "111110",      length => 6),
        (code => "1111110",     length => 7),
        (code => "11111110",    length => 8),
        (code => "111111110",   length => 9)
    );
    
    type ac_code_type is record
        code   : std_logic_vector(15 downto 0);
        length : integer range 0 to 16;
    end record;
    
    type ac_luma_array is array(0 to 15, 0 to 10) of ac_code_type;
    constant AC_LUMA_HUFF : ac_luma_array := (
    0 => (
        0 => (code => "1010", length => 4),
        1 => (code => "00", length => 2),
        2 => (code => "01", length => 2),
        3 => (code => "100", length => 3),
        4 => (code => "1011", length => 4),
        5 => (code => "11010", length => 5),
        6 => (code => "1111000", length => 7),
        7 => (code => "11111000", length => 8),
        8 => (code => "1111110110", length => 10),
        9 => (code => "1111111110000010", length => 16),
        10 => (code => "1111111110000011", length => 16),
        others => (code => (others => '0'), length => 0)  
    ),
    1 => (
        1 => (code => "1100", length => 4),
        2 => (code => "11011", length => 5),
        3 => (code => "1111001", length => 7),
        4 => (code => "111110110", length => 9),
        5 => (code => "11111110110", length => 11),
        6 => (code => "1111111110000100", length => 16),
        7 => (code => "1111111110000101", length => 16),
        8 => (code => "1111111110000110", length => 16),
        9 => (code => "1111111110000111", length => 16),
        10 => (code => "1111111110001000", length => 16),
        
        others => (code => (others => '0'), length => 0)
    ),
    2 => (
        1 => (code => "11100", length => 5),
        2 => (code => "11111001", length => 8),
        3 => (code => "1111110111", length => 10),
        4 => (code => "111111110100", length => 12),
        5 => (code => "1111111110001001", length => 16),
        6 => (code => "1111111110001010", length => 16),
        7 => (code => "1111111110001011", length => 16),
        8 => (code => "1111111110001100", length => 16),
        9 => (code => "1111111110001101", length => 16),
        10 => (code => "1111111110001110", length => 16),
        
        others => (code => (others => '0'), length => 0)
    ),
--        (3, 1):  ("111010",                6),
--        (3, 2):  ("111110111",             9),
--        (3, 3):  ("111111110101",         12),
--        (3, 4):  ("1111111110001111",      16),
--        (3, 5):  ("1111111110010000",      16),
--        (3, 6):  ("1111111110010001",      16),
--        (3, 7):  ("1111111110010010",      16),
--        (3, 8):  ("1111111110010011",      16),
--        (3, 9):  ("1111111110010100",      16),
--        (3, 10): ("1111111110010101",      16),
    
--        (4, 1):  ("111011",                6),
--        (4, 2):  ("1111111000",           10),
--        (4, 3):  ("1111111110010110",      16),
--        (4, 4):  ("1111111110010111",      16),
--        (4, 5):  ("1111111110011000",      16),
--        (4, 6):  ("1111111110011001",      16),
--        (4, 7):  ("1111111110011010",      16),
--        (4, 8):  ("1111111110011011",      16),
--        (4, 9):  ("1111111110011100",      16),
--        (4, 10): ("1111111110011101",      16),
    
--        (5, 1):  ("1111010",               7),
--        (5, 2):  ("11111110111",          11),
--        (5, 3):  ("1111111110011110",      16),
--        (5, 4):  ("1111111110011111",      16),
--        (5, 5):  ("1111111110100000",      16),
--        (5, 6):  ("1111111110100001",      16),
--        (5, 7):  ("1111111110100010",      16),
--        (5, 8):  ("1111111110100011",      16),
--        (5, 9):  ("1111111110100100",      16),
--        (5, 10): ("1111111110100101",      16),
    
--        (6, 1):  ("1111011",               7),
--        (6, 2):  ("111111110110",         12),
--        (6, 3):  ("1111111110100110",      16),
--        (6, 4):  ("1111111110100111",      16),
--        (6, 5):  ("1111111110101000",      16),
--        (6, 6):  ("1111111110101001",      16),
--        (6, 7):  ("1111111110101010",      16),
--        (6, 8):  ("1111111110101011",      16),
--        (6, 9):  ("1111111110101100",      16),
--        (6, 10): ("1111111110101101",      16),
    
--        (7, 1):  ("11111010",              8),
--        (7, 2):  ("111111110111",         12),
--        (7, 3):  ("1111111110101110",      16),
--        (7, 4):  ("1111111110101111",      16),
--        (7, 5):  ("1111111110110000",      16),
--        (7, 6):  ("1111111110110001",      16),
--        (7, 7):  ("1111111110110010",      16),
--        (7, 8):  ("1111111110110011",      16),
--        (7, 9):  ("1111111110110100",      16),
--        (7, 10): ("1111111110110101",      16),
    
--        (8, 1):  ("111111000",            10),
--        (8, 2):  ("111111111000000",      15),
--        (8, 3):  ("1111111110110110",      16),
--        (8, 4):  ("1111111110110111",      16),
--        (8, 5):  ("1111111110111000",      16),
--        (8, 6):  ("1111111110111001",      16),
--        (8, 7):  ("1111111110111010",      16),
--        (8, 8):  ("1111111110111011",      16),
--        (8, 9):  ("1111111110111100",      16),
--        (8, 10): ("1111111110111101",      16),
    
--        (9, 1):  ("111111001",            10),
--        (9, 2):  ("1111111110111110",      16),
--        (9, 3):  ("1111111110111111",      16),
--        (9, 4):  ("1111111111000000",      16),
--        (9, 5):  ("1111111111000001",      16),
--        (9, 6):  ("1111111111000010",      16),
--        (9, 7):  ("1111111111000011",      16),
--        (9, 8):  ("1111111111000100",      16),
--        (9, 9):  ("1111111111000101",      16),
--        (9, 10): ("1111111111000110",      16),
    
--        (10, 1): ("111111010",            10),
--        (10, 2): ("1111111111000111",      16),
--        (10, 3): ("1111111111001000",      16),
--        (10, 4): ("1111111111001001",      16),
--        (10, 5): ("1111111111001010",      16),
--        (10, 6): ("1111111111001011",      16),
--        (10, 7): ("1111111111001100",      16),
--        (10, 8): ("1111111111001101",      16),
--        (10, 9): ("1111111111001110",      16),
--        (10, 10):("1111111111001111",      16),
    
--        (11, 1): ("1111111001",           10),
--        (11, 2): ("1111111111010000",      16),
--        (11, 3): ("1111111111010001",      16),
--        (11, 4): ("1111111111010010",      16),
--        (11, 5): ("1111111111010011",      16),
--        (11, 6): ("1111111111010100",      16),
--        (11, 7): ("1111111111010101",      16),
--        (11, 8): ("1111111111010110",      16),
--        (11, 9): ("1111111111010111",      16),
--        (11, 10):("1111111111011000",      16),
    
--        (12, 1): ("1111111010",           10),
--        (12, 2): ("1111111111011001",      16),
--        (12, 3): ("1111111111011010",      16),
--        (12, 4): ("1111111111011011",      16),
--        (12, 5): ("1111111111011100",      16),
--        (12, 6): ("1111111111011101",      16),
--        (12, 7): ("1111111111011110",      16),
--        (12, 8): ("1111111111011111",      16),
--        (12, 9): ("1111111111100000",      16),
--        (12, 10):("1111111111100001",      16),
    
--        (13, 1): ("11111111000",          11),
--        (13, 2): ("1111111111100010",      16),
--        (13, 3): ("1111111111100011",      16),
--        (13, 4): ("1111111111100100",      16),
--        (13, 5): ("1111111111100101",      16),
--        (13, 6): ("1111111111100110",      16),
--        (13, 7): ("1111111111100111",      16),
--        (13, 8): ("1111111111101000",      16),
--        (13, 9): ("1111111111101001",      16),
--        (13, 10):("1111111111101010",      16),
    
--        (14, 1): ("1111111111101011",     16),
--        (14, 2): ("1111111111101100",      16),
--        (14, 3): ("1111111111101101",      16),
--        (14, 4): ("1111111111101110",      16),
--        (14, 5): ("1111111111101111",      16),
--        (14, 6): ("1111111111110000",      16),
--        (14, 7): ("1111111111110001",      16),
--        (14, 8): ("1111111111110010",      16),
--        (14, 9): ("1111111111110011",      16),
--        (14, 10):("1111111111110100",      16),
    
--        (15, 0): ("11111111001",          11),
--        (15, 1): ("1111111111110101",      16),
--        (15, 2): ("1111111111110110",      16),
--        (15, 3): ("1111111111110111",      16),
--        (15, 4): ("1111111111111000",      16),
--        (15, 5): ("1111111111111001",      16),
--        (15, 6): ("1111111111111010",      16),
--        (15, 7): ("1111111111111011",      16),
--        (15, 8): ("1111111111111100",      16),
--        (15, 9): ("1111111111111101",      16),
--        (15, 10):("1111111111111110",      16),


    );

end package;